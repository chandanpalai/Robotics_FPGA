----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    03:18:08 03/20/2013 
-- Design Name: 
-- Module Name:    compute_xy - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity compute_xy is
    Port ( done : in  STD_LOGIC;
           din : in  STD_LOGIC;
           i : in  STD_LOGIC;
           xin : in  STD_LOGIC;
           yin : in  STD_LOGIC;
           xout : in  STD_LOGIC;
           yout : in  STD_LOGIC;
           dout : in  STD_LOGIC;
           done : in  STD_LOGIC);
end compute_xy;

architecture Behavioral of compute_xy is

begin


end Behavioral;

